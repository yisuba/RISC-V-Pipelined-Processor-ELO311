
// Data_Memory
////// Solo Carcasa
////////////////////////////

module Data_Memory(
	input logic clk, rst, WE,
	input logic [31:0] A, WD,
	output logic [31:0] RD
);

endmodule