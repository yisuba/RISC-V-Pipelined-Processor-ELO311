`timescale 1ns / 1ps


///// 11/01/25
// Etapa de Execute 
////// 
////// 
////// 
////////////////////////////

module Execute_Stage(
	input logic [4:0] RD1E, RD2E, 
	input logic [4:0] Rs1E, Rs2E, RdE,
	input logic [2:0] ALUControlE,
	input logic [24:0] ExtImmE
	input logic [31:0] PCE, PCPlus4E
);
	
	

endmodule